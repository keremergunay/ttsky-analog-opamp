magic
tech sky130B
magscale 1 2
timestamp 1768741062
<< metal1 >>
rect 12240 32374 12250 32375
rect 12234 31981 12250 32374
rect 12644 31981 12654 32375
rect 12234 28558 12650 31981
rect 12245 27645 12640 28558
rect 43666 18051 43888 18052
rect 43664 17853 43674 18051
rect 43872 17853 43888 18051
rect 43666 16263 43888 17853
rect 14510 13082 15052 13092
rect 10156 13006 10852 13008
rect 10156 12996 11024 13006
rect 10156 12808 10916 12996
rect 11104 12808 11114 12996
rect 14510 12894 14944 13082
rect 15132 12894 15142 13082
rect 14510 12886 15052 12894
rect 10780 12800 11024 12808
rect 2850 4897 3054 6884
rect 2848 4711 2858 4897
rect 3044 4711 3054 4897
rect 2850 4710 3054 4711
rect 15074 1728 15287 2096
rect 15074 1515 15499 1728
rect 15286 1438 15499 1515
rect 14726 1426 15616 1438
rect 14726 1007 14742 1426
rect 15161 1007 15616 1426
rect 14726 990 15616 1007
<< via1 >>
rect 12250 31981 12644 32375
rect 43674 17853 43872 18051
rect 10916 12808 11104 12996
rect 14944 12894 15132 13082
rect 2858 4711 3044 4897
rect 14742 1007 15161 1426
<< metal2 >>
rect 12250 33002 12646 33012
rect 12250 32610 12254 33002
rect 12250 32600 12646 32610
rect 12250 32375 12644 32600
rect 12250 31971 12644 31981
rect 43682 18390 43870 18398
rect 43674 18388 43872 18390
rect 43674 18200 43682 18388
rect 43870 18200 43872 18388
rect 43674 18051 43872 18200
rect 43674 17843 43872 17853
rect 14944 13084 15132 13092
rect 15208 13084 15392 13086
rect 14944 13082 15394 13084
rect 10916 12998 11104 13006
rect 11180 12998 11364 13000
rect 10916 12996 11366 12998
rect 11104 12990 11366 12996
rect 11104 12808 11180 12990
rect 10916 12806 11180 12808
rect 11364 12806 11366 12990
rect 15132 13076 15394 13082
rect 15132 12894 15208 13076
rect 14944 12892 15208 12894
rect 15392 12892 15394 13076
rect 14944 12884 15132 12892
rect 15208 12882 15392 12892
rect 10916 12798 11104 12806
rect 11180 12796 11364 12806
rect 2858 4897 3044 4907
rect 2854 4711 2858 4734
rect 2854 4558 3044 4711
rect 2854 4548 3046 4558
rect 2854 4360 2858 4548
rect 2854 4358 3046 4360
rect 2858 4350 3046 4358
rect 14742 1426 15161 1436
rect 14325 1418 14742 1426
rect 13920 1408 14742 1418
rect 14336 1008 14742 1408
rect 14336 992 14350 1008
rect 14736 1007 14742 1008
rect 14742 997 15161 1007
rect 13920 990 14350 992
rect 13920 982 14336 990
<< via2 >>
rect 12254 32610 12646 33002
rect 43682 18200 43870 18388
rect 11180 12806 11364 12990
rect 15208 12892 15392 13076
rect 2858 4360 3046 4548
rect 13920 992 14336 1408
<< metal3 >>
rect 12254 33740 12646 33748
rect 12246 33340 12256 33740
rect 12656 33340 12666 33740
rect 12254 33007 12646 33340
rect 12244 33002 12656 33007
rect 12244 32610 12254 33002
rect 12646 32610 12656 33002
rect 12244 32605 12656 32610
rect 43682 18704 43870 18706
rect 43674 18524 43684 18704
rect 43864 18524 43874 18704
rect 43682 18393 43870 18524
rect 43672 18388 43880 18393
rect 43672 18200 43682 18388
rect 43870 18200 43880 18388
rect 43672 18195 43880 18200
rect 15198 13076 15402 13081
rect 11170 12990 11374 12995
rect 11170 12806 11180 12990
rect 11364 12810 11476 12990
rect 11656 12810 11666 12990
rect 15198 12892 15208 13076
rect 15392 12896 15504 13076
rect 15684 12896 15694 13076
rect 15392 12892 15684 12896
rect 15198 12887 15402 12892
rect 11364 12806 11656 12810
rect 11170 12801 11374 12806
rect 2848 4548 3056 4553
rect 2848 4360 2858 4548
rect 3046 4360 3056 4548
rect 2848 4355 3056 4360
rect 2858 4236 3046 4355
rect 2844 4056 2854 4236
rect 3034 4056 3046 4236
rect 2858 4048 3046 4056
rect 13910 1408 14346 1413
rect 13220 1400 13920 1408
rect 13220 1000 13240 1400
rect 13640 1000 13920 1400
rect 13220 992 13920 1000
rect 14336 992 14346 1408
rect 13220 987 14346 992
rect 13220 978 14056 987
<< via3 >>
rect 12256 33340 12656 33740
rect 43684 18524 43864 18704
rect 11476 12810 11656 12990
rect 15504 12896 15684 13076
rect 2854 4056 3034 4236
rect 13240 1000 13640 1400
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 44384 4786 44784
rect 200 1000 600 44384
rect 800 1400 1200 44152
rect 4386 34594 4786 44384
rect 4386 34194 12656 34594
rect 12256 33741 12656 34194
rect 12255 33740 12657 33741
rect 12255 33340 12256 33740
rect 12656 33340 12657 33740
rect 12255 33339 12657 33340
rect 6800 26994 40628 27174
rect 6800 8522 6980 26994
rect 40448 23054 40628 26994
rect 40448 22874 41044 23054
rect 40864 18704 41044 22874
rect 43683 18704 43865 18705
rect 40864 18524 43684 18704
rect 43864 18524 43865 18704
rect 43683 18523 43865 18524
rect 15503 13076 15685 13077
rect 11646 12991 12776 13000
rect 11475 12990 12776 12991
rect 11475 12810 11476 12990
rect 11656 12820 12776 12990
rect 15503 12896 15504 13076
rect 15684 12896 25246 13076
rect 15503 12895 15685 12896
rect 11656 12810 11770 12820
rect 11475 12809 11657 12810
rect 12596 11060 12776 12820
rect 12596 10880 23938 11060
rect 6800 8342 17624 8522
rect 2853 4236 3035 4237
rect 2853 4056 2854 4236
rect 3034 4056 3035 4236
rect 2853 4055 3035 4056
rect 2854 3992 3034 4055
rect 2854 3812 16766 3992
rect 13239 1400 13641 1401
rect 800 1000 13240 1400
rect 13640 1000 13641 1400
rect 13239 999 13641 1000
rect 16586 668 16766 3812
rect 17444 2552 17624 8342
rect 23758 7910 23938 10880
rect 25066 8680 25246 12896
rect 25066 8500 30542 8680
rect 23758 7730 26678 7910
rect 17444 2372 22814 2552
rect 16586 488 18950 668
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 488
rect 22634 0 22814 2372
rect 26498 0 26678 7730
rect 30362 0 30542 8500
use two_stage_opamp  two_stage_opamp_0 Final_Project
timestamp 1768091639
transform 1 0 -306 0 1 11038
box 3266 -9126 44228 16662
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 1000 600 44152 1 FreeSans 2 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1768749653
<< metal1 >>
rect 12040 32374 12050 32375
rect 12034 31981 12050 32374
rect 12444 31981 12454 32375
rect 12034 28558 12450 31981
rect 12045 27645 12440 28558
rect 43466 18051 43688 18052
rect 43464 17853 43474 18051
rect 43672 17853 43688 18051
rect 43466 16263 43688 17853
rect 14310 13082 14852 13092
rect 9956 13006 10652 13008
rect 9956 12996 10824 13006
rect 9956 12808 10716 12996
rect 10904 12808 10914 12996
rect 14310 12894 14744 13082
rect 14932 12894 14942 13082
rect 14310 12886 14852 12894
rect 10580 12800 10824 12808
rect 2650 6680 3146 6884
rect 2650 4897 2854 6680
rect 2648 4711 2658 4897
rect 2844 4711 2854 4897
rect 2650 4710 2854 4711
rect 14874 1728 15087 2096
rect 14874 1515 15299 1728
rect 15086 1438 15299 1515
rect 14526 1426 15416 1438
rect 14526 1007 14542 1426
rect 14961 1007 15416 1426
rect 14526 990 15416 1007
<< via1 >>
rect 12050 31981 12444 32375
rect 43474 17853 43672 18051
rect 10716 12808 10904 12996
rect 14744 12894 14932 13082
rect 2658 4711 2844 4897
rect 14542 1007 14961 1426
<< metal2 >>
rect 12050 33002 12446 33012
rect 12050 32610 12054 33002
rect 12050 32600 12446 32610
rect 12050 32375 12444 32600
rect 12050 31971 12444 31981
rect 43482 18390 43670 18398
rect 43474 18388 43672 18390
rect 43474 18200 43482 18388
rect 43670 18200 43672 18388
rect 43474 18051 43672 18200
rect 43474 17843 43672 17853
rect 14744 13084 14932 13092
rect 15008 13084 15192 13086
rect 14744 13082 15194 13084
rect 10716 12998 10904 13006
rect 10980 12998 11164 13000
rect 10716 12996 11166 12998
rect 10904 12990 11166 12996
rect 10904 12808 10980 12990
rect 10716 12806 10980 12808
rect 11164 12806 11166 12990
rect 14932 13076 15194 13082
rect 14932 12894 15008 13076
rect 14744 12892 15008 12894
rect 15192 12892 15194 13076
rect 14744 12884 14932 12892
rect 15008 12882 15192 12892
rect 10716 12798 10904 12806
rect 10980 12796 11164 12806
rect 2658 4897 2844 4907
rect 2654 4711 2658 4734
rect 2654 4558 2844 4711
rect 2654 4548 2846 4558
rect 2654 4360 2658 4548
rect 2654 4358 2846 4360
rect 2658 4350 2846 4358
rect 14542 1426 14961 1436
rect 14125 1418 14542 1426
rect 13720 1408 14542 1418
rect 14136 1008 14542 1408
rect 14136 992 14150 1008
rect 14536 1007 14542 1008
rect 14542 997 14961 1007
rect 13720 990 14150 992
rect 13720 982 14136 990
<< via2 >>
rect 12054 32610 12446 33002
rect 43482 18200 43670 18388
rect 10980 12806 11164 12990
rect 15008 12892 15192 13076
rect 2658 4360 2846 4548
rect 13720 992 14136 1408
<< metal3 >>
rect 12054 33740 12446 33748
rect 12046 33340 12056 33740
rect 12456 33340 12466 33740
rect 12054 33007 12446 33340
rect 12044 33002 12456 33007
rect 12044 32610 12054 33002
rect 12446 32610 12456 33002
rect 12044 32605 12456 32610
rect 43482 18704 43670 18706
rect 43474 18524 43484 18704
rect 43664 18524 43674 18704
rect 43482 18393 43670 18524
rect 43472 18388 43680 18393
rect 43472 18200 43482 18388
rect 43670 18200 43680 18388
rect 43472 18195 43680 18200
rect 14998 13076 15202 13081
rect 10970 12990 11174 12995
rect 10970 12806 10980 12990
rect 11164 12810 11276 12990
rect 11456 12810 11466 12990
rect 14998 12892 15008 13076
rect 15192 12896 15304 13076
rect 15484 12896 15494 13076
rect 15192 12892 15484 12896
rect 14998 12887 15202 12892
rect 11164 12806 11456 12810
rect 10970 12801 11174 12806
rect 2648 4548 2856 4553
rect 2648 4360 2658 4548
rect 2846 4360 2856 4548
rect 2648 4355 2856 4360
rect 2658 4236 2846 4355
rect 2644 4056 2654 4236
rect 2834 4056 2846 4236
rect 2658 4048 2846 4056
rect 13710 1408 14146 1413
rect 13020 1400 13720 1408
rect 13020 1000 13040 1400
rect 13440 1000 13720 1400
rect 13020 992 13720 1000
rect 14136 992 14146 1408
rect 13020 987 14146 992
rect 13020 978 13856 987
<< via3 >>
rect 12056 33340 12456 33740
rect 43484 18524 43664 18704
rect 11276 12810 11456 12990
rect 15304 12896 15484 13076
rect 2654 4056 2834 4236
rect 13040 1000 13440 1400
<< metal4 >>
rect 5934 44952 5994 45152
rect 6486 44952 6546 45152
rect 7038 44952 7098 45152
rect 7590 44952 7650 45152
rect 8142 44952 8202 45152
rect 8694 44952 8754 45152
rect 9246 44952 9306 45152
rect 9798 44952 9858 45152
rect 10350 44952 10410 45152
rect 10902 44952 10962 45152
rect 11454 44952 11514 45152
rect 12006 44952 12066 45152
rect 12558 44952 12618 45152
rect 13110 44952 13170 45152
rect 13662 44952 13722 45152
rect 14214 44952 14274 45152
rect 14766 44952 14826 45152
rect 15318 44952 15378 45152
rect 15870 44952 15930 45152
rect 16422 44952 16482 45152
rect 16974 44952 17034 45152
rect 17526 44952 17586 45152
rect 18078 44952 18138 45152
rect 18630 44952 18690 45152
rect 19182 44952 19242 45152
rect 19734 44952 19794 45152
rect 20286 44952 20346 45152
rect 20838 44952 20898 45152
rect 21390 44952 21450 45152
rect 21942 44952 22002 45152
rect 22494 44952 22554 45152
rect 23046 44952 23106 45152
rect 23598 44952 23658 45152
rect 24150 44952 24210 45152
rect 24702 44952 24762 45152
rect 25254 44952 25314 45152
rect 25806 44952 25866 45152
rect 26358 44952 26418 45152
rect 26910 44952 26970 45152
rect 27462 44952 27522 45152
rect 28014 44952 28074 45152
rect 28566 44952 28626 45152
rect 29118 44952 29178 45152
rect 0 44384 4586 44784
rect 0 1000 400 44384
rect 600 1400 1000 44152
rect 4186 34594 4586 44384
rect 4186 34194 12456 34594
rect 12056 33741 12456 34194
rect 12055 33740 12457 33741
rect 12055 33340 12056 33740
rect 12456 33340 12457 33740
rect 12055 33339 12457 33340
rect 6600 26994 40428 27174
rect 6600 8522 6780 26994
rect 40248 23054 40428 26994
rect 40248 22874 40844 23054
rect 40664 18704 40844 22874
rect 43483 18704 43665 18705
rect 40664 18524 43484 18704
rect 43664 18524 43665 18704
rect 43483 18523 43665 18524
rect 15303 13076 15485 13077
rect 11446 12991 12576 13000
rect 11275 12990 12576 12991
rect 11275 12810 11276 12990
rect 11456 12820 12576 12990
rect 15303 12896 15304 13076
rect 15484 12896 25046 13076
rect 15303 12895 15485 12896
rect 11456 12810 11570 12820
rect 11275 12809 11457 12810
rect 12396 11060 12576 12820
rect 12396 10880 23738 11060
rect 6600 8342 17424 8522
rect 2653 4236 2835 4237
rect 2653 4056 2654 4236
rect 2834 4056 2835 4236
rect 2653 4055 2835 4056
rect 2654 3992 2834 4055
rect 2654 3812 16566 3992
rect 13039 1400 13441 1401
rect 600 1000 13040 1400
rect 13440 1000 13441 1400
rect 13039 999 13441 1000
rect 16386 668 16566 3812
rect 17244 2552 17424 8342
rect 23558 7910 23738 10880
rect 24866 8680 25046 12896
rect 24866 8500 30342 8680
rect 23558 7730 26478 7910
rect 17244 2372 22614 2552
rect 16386 488 18750 668
rect 3114 0 3294 200
rect 6978 0 7158 200
rect 10842 0 11022 200
rect 14706 0 14886 200
rect 18570 0 18750 488
rect 22434 0 22614 2372
rect 26298 0 26478 7730
rect 30162 0 30342 8500
use two_stage_opamp  two_stage_opamp_0 ~/Desktop/design/mag/Final_Project
timestamp 1768091639
transform 1 0 -306 0 1 11036
box 3266 -9126 44228 16662
<< labels >>
flabel metal4 s 28566 44952 28626 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29118 44952 29178 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28014 44952 28074 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30162 0 30342 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26298 0 26478 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22434 0 22614 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18570 0 18750 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14706 0 14886 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 10842 0 11022 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 6978 0 7158 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3114 0 3294 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27462 44952 27522 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 26910 44952 26970 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26358 44952 26418 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 25806 44952 25866 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25254 44952 25314 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24702 44952 24762 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24150 44952 24210 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23598 44952 23658 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23046 44952 23106 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22494 44952 22554 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 21942 44952 22002 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21390 44952 21450 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20838 44952 20898 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20286 44952 20346 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19734 44952 19794 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19182 44952 19242 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9798 44952 9858 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 9246 44952 9306 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 8694 44952 8754 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 8142 44952 8202 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 7590 44952 7650 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 7038 44952 7098 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 6486 44952 6546 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 5934 44952 5994 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 14214 44952 14274 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 13662 44952 13722 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 13110 44952 13170 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 12558 44952 12618 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 12006 44952 12066 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 11454 44952 11514 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 10902 44952 10962 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 10350 44952 10410 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 18630 44952 18690 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 18078 44952 18138 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 17526 44952 17586 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 16974 44952 17034 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 16422 44952 16482 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 15870 44952 15930 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 15318 44952 15378 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 14766 44952 14826 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 0 1000 400 44152 1 FreeSans 2 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 600 1000 1000 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>

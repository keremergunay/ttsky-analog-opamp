VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_keremergunay_two_stage_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_keremergunay_two_stage_opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 334.880 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 142.830 224.760 143.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 145.590 224.760 145.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.070 224.760 140.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER li1 ;
        RECT 72.590 63.030 73.590 63.200 ;
      LAYER mcon ;
        RECT 72.670 63.030 73.510 63.200 ;
      LAYER met1 ;
        RECT 71.550 65.410 74.260 65.460 ;
        RECT 71.550 64.470 74.710 65.410 ;
        RECT 71.550 64.430 74.260 64.470 ;
        RECT 72.560 63.970 73.560 64.430 ;
        RECT 72.940 63.230 73.260 63.970 ;
        RECT 72.610 63.000 73.570 63.230 ;
      LAYER via ;
        RECT 73.720 64.470 74.660 65.410 ;
      LAYER met2 ;
        RECT 73.720 65.420 74.660 65.460 ;
        RECT 75.040 65.420 75.960 65.430 ;
        RECT 73.720 64.460 75.970 65.420 ;
        RECT 73.720 64.420 74.660 64.460 ;
        RECT 75.040 64.410 75.960 64.460 ;
      LAYER via2 ;
        RECT 75.040 64.460 75.960 65.380 ;
      LAYER met3 ;
        RECT 74.990 65.380 76.010 65.405 ;
        RECT 74.990 64.480 77.470 65.380 ;
        RECT 74.990 64.460 77.420 64.480 ;
        RECT 74.990 64.435 76.010 64.460 ;
      LAYER via3 ;
        RECT 76.520 64.480 77.420 65.380 ;
      LAYER met4 ;
        RECT 76.515 65.380 77.425 65.385 ;
        RECT 76.515 64.480 125.230 65.380 ;
        RECT 76.515 64.475 77.425 64.480 ;
        RECT 124.330 43.400 125.230 64.480 ;
        RECT 124.330 42.500 151.710 43.400 ;
        RECT 150.810 0.000 151.710 42.500 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER li1 ;
        RECT 50.800 62.990 51.800 63.160 ;
      LAYER mcon ;
        RECT 50.880 62.990 51.720 63.160 ;
      LAYER met1 ;
        RECT 49.780 65.030 53.260 65.040 ;
        RECT 49.780 64.980 54.120 65.030 ;
        RECT 49.780 64.040 54.570 64.980 ;
        RECT 50.780 64.030 51.780 64.040 ;
        RECT 51.160 63.190 51.440 64.030 ;
        RECT 52.900 64.000 54.120 64.040 ;
        RECT 50.820 62.960 51.780 63.190 ;
      LAYER via ;
        RECT 53.580 64.040 54.520 64.980 ;
      LAYER met2 ;
        RECT 53.580 64.990 54.520 65.030 ;
        RECT 54.900 64.990 55.820 65.000 ;
        RECT 53.580 64.030 55.830 64.990 ;
        RECT 53.580 63.990 54.520 64.030 ;
        RECT 54.900 63.980 55.820 64.030 ;
      LAYER via2 ;
        RECT 54.900 64.030 55.820 64.950 ;
      LAYER met3 ;
        RECT 54.850 64.950 55.870 64.975 ;
        RECT 54.850 64.050 57.330 64.950 ;
        RECT 54.850 64.030 57.280 64.050 ;
        RECT 54.850 64.005 55.870 64.030 ;
      LAYER via3 ;
        RECT 56.380 64.050 57.280 64.950 ;
      LAYER met4 ;
        RECT 57.230 64.955 62.880 65.000 ;
        RECT 56.375 64.100 62.880 64.955 ;
        RECT 56.375 64.050 57.850 64.100 ;
        RECT 56.375 64.045 57.285 64.050 ;
        RECT 61.980 55.300 62.880 64.100 ;
        RECT 61.980 54.400 118.690 55.300 ;
        RECT 117.790 39.550 118.690 54.400 ;
        RECT 117.790 38.650 132.390 39.550 ;
        RECT 131.490 0.000 132.390 38.650 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.710199 ;
    PORT
      LAYER li1 ;
        RECT 209.440 110.790 209.610 135.210 ;
        RECT 207.090 17.390 207.260 33.430 ;
      LAYER mcon ;
        RECT 209.440 110.870 209.610 135.130 ;
        RECT 207.090 17.470 207.260 33.350 ;
      LAYER met1 ;
        RECT 209.410 120.405 209.640 135.190 ;
        RECT 197.315 118.555 209.640 120.405 ;
        RECT 197.315 83.540 199.165 118.555 ;
        RECT 209.410 110.810 209.640 118.555 ;
        RECT 217.330 90.255 218.440 90.260 ;
        RECT 217.320 89.265 218.440 90.255 ;
        RECT 197.315 83.110 203.370 83.540 ;
        RECT 192.480 82.560 203.370 83.110 ;
        RECT 192.480 81.260 199.165 82.560 ;
        RECT 202.390 82.230 203.370 82.560 ;
        RECT 217.330 82.230 218.440 89.265 ;
        RECT 218.610 82.230 219.610 82.270 ;
        RECT 202.390 81.270 219.610 82.230 ;
        RECT 192.540 81.210 194.540 81.260 ;
        RECT 202.390 81.250 219.040 81.270 ;
        RECT 202.390 35.600 203.370 81.250 ;
        RECT 202.340 34.640 203.400 35.600 ;
        RECT 202.390 34.630 203.370 34.640 ;
        RECT 202.345 28.925 203.375 29.855 ;
        RECT 202.395 25.520 203.325 28.925 ;
        RECT 207.060 25.520 207.290 33.410 ;
        RECT 202.395 24.590 207.290 25.520 ;
        RECT 207.060 17.410 207.290 24.590 ;
      LAYER via ;
        RECT 217.370 89.265 218.360 90.255 ;
        RECT 192.590 81.210 194.490 83.110 ;
        RECT 202.390 34.640 203.350 35.600 ;
        RECT 202.395 28.925 203.325 29.855 ;
      LAYER met2 ;
        RECT 217.410 91.950 218.350 91.990 ;
        RECT 217.370 89.215 218.360 91.950 ;
        RECT 189.110 83.110 190.960 83.160 ;
        RECT 192.590 83.110 194.490 83.160 ;
        RECT 189.060 81.210 194.490 83.110 ;
        RECT 192.590 81.160 194.490 81.210 ;
        RECT 202.390 29.860 203.350 35.650 ;
        RECT 202.390 28.910 203.340 29.860 ;
        RECT 202.395 28.875 203.325 28.910 ;
      LAYER via2 ;
        RECT 217.410 91.000 218.350 91.940 ;
        RECT 189.110 81.260 190.960 83.110 ;
      LAYER met3 ;
        RECT 131.700 116.040 185.950 116.210 ;
        RECT 131.700 115.610 186.085 116.040 ;
        RECT 131.700 85.320 158.085 115.610 ;
        RECT 131.870 85.040 158.085 85.320 ;
        RECT 159.930 85.040 186.085 115.610 ;
        RECT 217.410 93.520 218.350 93.530 ;
        RECT 217.370 92.620 218.370 93.520 ;
        RECT 217.410 91.965 218.350 92.620 ;
        RECT 217.360 90.975 218.400 91.965 ;
        RECT 131.870 78.040 132.470 85.040 ;
        RECT 185.350 83.110 185.950 85.040 ;
        RECT 189.060 83.110 191.010 83.135 ;
        RECT 185.300 81.260 191.010 83.110 ;
        RECT 185.350 78.040 185.950 81.260 ;
        RECT 189.060 81.235 191.010 81.260 ;
        RECT 131.870 47.470 158.085 78.040 ;
        RECT 159.930 47.470 186.085 78.040 ;
        RECT 131.870 47.040 186.085 47.470 ;
        RECT 131.870 46.870 186.070 47.040 ;
      LAYER via3 ;
        RECT 157.665 85.180 157.985 115.900 ;
        RECT 185.665 85.180 185.985 115.900 ;
        RECT 217.420 92.620 218.320 93.520 ;
        RECT 157.665 47.180 157.985 77.900 ;
        RECT 185.665 47.180 185.985 77.900 ;
      LAYER met4 ;
        RECT 33.000 134.970 202.140 135.870 ;
        RECT 33.000 42.610 33.900 134.970 ;
        RECT 157.585 85.100 158.065 115.980 ;
        RECT 185.585 85.100 186.065 115.980 ;
        RECT 201.240 115.270 202.140 134.970 ;
        RECT 201.240 114.370 204.220 115.270 ;
        RECT 203.320 93.520 204.220 114.370 ;
        RECT 217.415 93.520 218.325 93.525 ;
        RECT 203.320 92.620 218.325 93.520 ;
        RECT 217.415 92.615 218.325 92.620 ;
        RECT 157.585 47.100 158.065 77.980 ;
        RECT 185.585 47.100 186.065 77.980 ;
        RECT 33.000 41.710 87.120 42.610 ;
        RECT 86.220 12.760 87.120 41.710 ;
        RECT 86.220 11.860 113.070 12.760 ;
        RECT 112.170 0.000 113.070 11.860 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 29.000000 ;
    ANTENNADIFFAREA 1.740000 ;
    PORT
      LAYER li1 ;
        RECT 26.445 41.390 26.615 41.890 ;
        RECT 24.190 41.160 26.230 41.330 ;
        RECT 18.025 33.545 18.525 33.715 ;
        RECT 32.235 33.475 32.735 33.645 ;
        RECT 61.040 33.570 61.540 33.740 ;
        RECT 110.920 33.570 111.420 33.740 ;
        RECT 207.320 33.600 208.320 33.770 ;
        RECT 17.795 31.335 17.965 33.375 ;
        RECT 32.005 31.265 32.175 33.305 ;
      LAYER mcon ;
        RECT 26.445 41.470 26.615 41.810 ;
        RECT 24.270 41.160 26.150 41.330 ;
        RECT 18.105 33.545 18.445 33.715 ;
        RECT 32.315 33.475 32.655 33.645 ;
        RECT 61.120 33.570 61.460 33.740 ;
        RECT 111.000 33.570 111.340 33.740 ;
        RECT 207.400 33.600 208.240 33.770 ;
        RECT 17.795 31.415 17.965 33.295 ;
        RECT 32.005 31.345 32.175 33.225 ;
      LAYER met1 ;
        RECT 26.415 41.780 26.645 41.870 ;
        RECT 26.415 41.410 26.720 41.780 ;
        RECT 24.210 41.130 26.210 41.360 ;
        RECT 24.950 39.810 25.190 41.130 ;
        RECT 26.480 39.810 26.720 41.410 ;
        RECT 24.950 39.570 26.720 39.810 ;
        RECT 13.250 34.380 15.730 34.420 ;
        RECT 13.250 33.800 15.800 34.380 ;
        RECT 24.950 33.800 25.190 39.570 ;
        RECT 13.250 33.570 208.300 33.800 ;
        RECT 13.250 33.560 208.270 33.570 ;
        RECT 13.250 33.400 15.800 33.560 ;
        RECT 13.250 24.485 14.270 33.400 ;
        RECT 14.800 33.380 15.800 33.400 ;
        RECT 16.630 32.540 16.900 33.560 ;
        RECT 18.045 33.515 18.505 33.560 ;
        RECT 17.765 32.540 17.995 33.355 ;
        RECT 16.630 32.270 17.995 32.540 ;
        RECT 30.470 32.640 30.710 33.560 ;
        RECT 32.255 33.445 32.715 33.560 ;
        RECT 61.060 33.540 61.520 33.560 ;
        RECT 110.940 33.540 111.400 33.560 ;
        RECT 31.975 32.640 32.205 33.285 ;
        RECT 30.470 32.400 32.205 32.640 ;
        RECT 17.765 31.355 17.995 32.270 ;
        RECT 31.975 31.285 32.205 32.400 ;
        RECT 13.240 23.555 14.270 24.485 ;
        RECT 13.250 23.550 14.270 23.555 ;
      LAYER via ;
        RECT 13.290 23.555 14.220 24.485 ;
      LAYER met2 ;
        RECT 13.290 23.670 14.220 24.535 ;
        RECT 13.270 22.790 14.220 23.670 ;
        RECT 13.270 21.790 14.230 22.790 ;
        RECT 13.290 21.750 14.230 21.790 ;
      LAYER via2 ;
        RECT 13.290 21.800 14.230 22.740 ;
      LAYER met3 ;
        RECT 13.240 21.775 14.280 22.765 ;
        RECT 13.290 21.180 14.230 21.775 ;
        RECT 13.220 20.280 14.230 21.180 ;
        RECT 13.290 20.240 14.230 20.280 ;
      LAYER via3 ;
        RECT 13.270 20.280 14.170 21.180 ;
      LAYER met4 ;
        RECT 13.265 20.275 14.175 21.185 ;
        RECT 13.270 19.960 14.170 20.275 ;
        RECT 13.270 19.060 82.830 19.960 ;
        RECT 81.930 3.340 82.830 19.060 ;
        RECT 81.930 2.440 93.750 3.340 ;
        RECT 92.850 0.000 93.750 2.440 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.530 0.000 74.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.210 0.000 55.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.890 0.000 35.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.570 0.000 16.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 137.310 224.760 137.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.550 224.760 134.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 131.790 224.760 132.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.030 224.760 129.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 126.270 224.760 126.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 123.510 224.760 123.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 120.750 224.760 121.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.990 224.760 118.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.230 224.760 115.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.470 224.760 112.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.710 224.760 110.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.950 224.760 107.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.190 224.760 104.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.430 224.760 101.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.670 224.760 98.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.910 224.760 96.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.990 224.760 49.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.230 224.760 46.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 43.470 224.760 43.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.710 224.760 41.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.950 224.760 38.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.190 224.760 35.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.430 224.760 32.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.670 224.760 29.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 71.070 224.760 71.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.310 224.760 68.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 65.550 224.760 65.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.790 224.760 63.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 60.030 224.760 60.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 57.270 224.760 57.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.510 224.760 54.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.750 224.760 52.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.150 224.760 93.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.390 224.760 90.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.630 224.760 87.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.870 224.760 85.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 82.110 224.760 82.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 79.350 224.760 79.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 76.590 224.760 76.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.830 224.760 74.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 221.920 22.930 223.920 ;
        RECT 0.000 5.000 2.000 221.920 ;
        RECT 20.930 172.970 22.930 221.920 ;
        RECT 20.930 170.970 62.280 172.970 ;
        RECT 60.280 168.705 62.280 170.970 ;
        RECT 60.275 166.695 62.285 168.705 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.000 7.000 5.000 220.760 ;
        RECT 65.195 7.000 67.205 7.005 ;
        RECT 3.000 5.000 67.205 7.000 ;
        RECT 65.195 4.995 67.205 5.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 48.650 71.560 48.820 131.600 ;
        RECT 70.230 71.530 70.400 131.570 ;
        RECT 90.720 112.430 90.890 117.470 ;
        RECT 90.950 112.045 91.450 112.215 ;
        RECT 209.670 110.405 210.170 110.575 ;
        RECT 115.095 84.890 115.425 85.060 ;
        RECT 114.930 79.680 115.100 84.720 ;
        RECT 115.420 79.680 115.590 84.720 ;
        RECT 48.880 71.175 53.880 71.345 ;
        RECT 70.460 71.145 75.460 71.315 ;
        RECT 50.570 59.780 50.740 62.820 ;
        RECT 51.860 59.780 52.030 62.820 ;
        RECT 72.360 59.820 72.530 62.860 ;
        RECT 73.650 59.820 73.820 62.860 ;
        RECT 26.445 54.100 26.615 54.600 ;
        RECT 24.190 53.870 26.230 54.040 ;
        RECT 24.120 48.530 26.160 48.700 ;
        RECT 26.375 47.970 26.545 48.470 ;
        RECT 24.120 47.740 26.160 47.910 ;
        RECT 24.190 41.950 26.230 42.120 ;
        RECT 60.810 29.360 60.980 33.400 ;
        RECT 110.690 17.360 110.860 33.400 ;
      LAYER mcon ;
        RECT 48.650 71.640 48.820 131.520 ;
        RECT 70.230 71.610 70.400 131.490 ;
        RECT 90.720 112.510 90.890 117.390 ;
        RECT 91.030 112.045 91.370 112.215 ;
        RECT 209.750 110.405 210.090 110.575 ;
        RECT 115.175 84.890 115.345 85.060 ;
        RECT 114.930 79.760 115.100 84.640 ;
        RECT 115.420 79.760 115.590 84.640 ;
        RECT 48.960 71.175 53.800 71.345 ;
        RECT 70.540 71.145 75.380 71.315 ;
        RECT 50.570 59.860 50.740 62.740 ;
        RECT 51.860 59.860 52.030 62.740 ;
        RECT 72.360 59.900 72.530 62.780 ;
        RECT 73.650 59.900 73.820 62.780 ;
        RECT 26.445 54.180 26.615 54.520 ;
        RECT 24.270 53.870 26.150 54.040 ;
        RECT 24.200 48.530 26.080 48.700 ;
        RECT 26.375 48.050 26.545 48.390 ;
        RECT 24.200 47.740 26.080 47.910 ;
        RECT 24.270 41.950 26.150 42.120 ;
        RECT 60.810 29.440 60.980 33.320 ;
        RECT 110.690 17.440 110.860 33.320 ;
      LAYER met1 ;
        RECT 48.620 82.720 48.850 131.580 ;
        RECT 43.150 82.220 48.850 82.720 ;
        RECT 43.150 68.190 43.650 82.220 ;
        RECT 48.620 71.580 48.850 82.220 ;
        RECT 70.200 74.265 70.430 131.550 ;
        RECT 101.260 120.855 190.875 121.200 ;
        RECT 90.690 114.600 90.920 117.450 ;
        RECT 65.930 73.695 70.430 74.265 ;
        RECT 48.900 71.145 53.860 71.375 ;
        RECT 50.960 68.190 51.460 71.145 ;
        RECT 65.930 70.200 66.500 73.695 ;
        RECT 70.200 71.550 70.430 73.695 ;
        RECT 81.780 113.640 90.920 114.600 ;
        RECT 70.480 71.115 75.440 71.345 ;
        RECT 65.890 69.660 66.530 70.200 ;
        RECT 72.780 68.190 73.280 71.115 ;
        RECT 81.780 70.565 82.740 113.640 ;
        RECT 90.690 112.450 90.920 113.640 ;
        RECT 90.970 112.190 91.430 112.245 ;
        RECT 90.970 112.015 91.480 112.190 ;
        RECT 90.980 103.170 91.480 112.015 ;
        RECT 85.870 102.670 91.480 103.170 ;
        RECT 81.740 69.615 82.790 70.565 ;
        RECT 81.780 69.600 82.740 69.615 ;
        RECT 85.870 68.190 86.370 102.670 ;
        RECT 101.260 95.235 101.605 120.855 ;
        RECT 190.530 109.490 190.875 120.855 ;
        RECT 209.690 110.375 210.150 110.605 ;
        RECT 209.730 109.520 210.130 110.375 ;
        RECT 195.360 109.490 196.165 109.520 ;
        RECT 190.530 109.145 196.165 109.490 ;
        RECT 195.360 109.110 196.165 109.145 ;
        RECT 202.070 109.120 210.130 109.520 ;
        RECT 195.360 109.100 196.120 109.110 ;
        RECT 43.150 67.690 86.370 68.190 ;
        RECT 90.730 94.890 101.605 95.235 ;
        RECT 43.150 61.300 43.650 67.690 ;
        RECT 69.705 66.035 79.600 66.425 ;
        RECT 65.900 63.860 66.540 64.400 ;
        RECT 50.540 61.300 50.770 62.800 ;
        RECT 43.150 60.800 50.770 61.300 ;
        RECT 50.540 59.800 50.770 60.800 ;
        RECT 51.830 61.270 52.060 62.800 ;
        RECT 65.950 61.440 66.490 63.860 ;
        RECT 69.705 61.440 70.095 66.035 ;
        RECT 72.330 61.440 72.560 62.840 ;
        RECT 51.830 60.910 59.330 61.270 ;
        RECT 51.830 59.800 52.060 60.910 ;
        RECT 24.210 53.840 26.210 54.070 ;
        RECT 24.950 52.670 25.250 53.840 ;
        RECT 26.390 52.670 26.690 54.630 ;
        RECT 24.950 52.370 26.690 52.670 ;
        RECT 24.950 48.730 25.250 52.370 ;
        RECT 58.970 51.820 59.330 60.910 ;
        RECT 65.950 60.900 72.560 61.440 ;
        RECT 72.330 59.840 72.560 60.900 ;
        RECT 73.620 61.440 73.850 62.840 ;
        RECT 73.620 61.080 77.070 61.440 ;
        RECT 73.620 59.840 73.850 61.080 ;
        RECT 76.710 51.820 77.070 61.080 ;
        RECT 79.210 56.940 79.600 66.035 ;
        RECT 81.760 61.770 82.780 62.690 ;
        RECT 79.210 56.930 80.190 56.940 ;
        RECT 79.210 56.560 80.235 56.930 ;
        RECT 79.210 56.550 80.190 56.560 ;
        RECT 58.970 51.460 77.070 51.820 ;
        RECT 24.140 48.500 26.140 48.730 ;
        RECT 26.345 48.430 26.575 48.450 ;
        RECT 26.345 47.990 26.700 48.430 ;
        RECT 24.140 47.710 26.140 47.940 ;
        RECT 24.950 45.550 25.210 47.710 ;
        RECT 26.440 45.550 26.700 47.990 ;
        RECT 24.950 45.290 45.160 45.550 ;
        RECT 48.830 45.290 57.370 45.550 ;
        RECT 24.950 42.150 25.210 45.290 ;
        RECT 24.210 41.920 26.210 42.150 ;
        RECT 58.970 35.660 59.330 51.460 ;
        RECT 60.215 45.265 77.725 45.570 ;
        RECT 60.270 45.260 77.725 45.265 ;
        RECT 81.810 38.590 82.730 61.770 ;
        RECT 90.730 56.925 91.075 94.890 ;
        RECT 85.270 56.580 91.075 56.925 ;
        RECT 96.940 86.760 115.360 87.080 ;
        RECT 96.940 45.570 97.260 86.760 ;
        RECT 115.040 85.090 115.360 86.760 ;
        RECT 115.040 84.860 115.405 85.090 ;
        RECT 115.040 84.840 115.360 84.860 ;
        RECT 114.900 80.770 115.130 84.700 ;
        RECT 83.980 45.250 97.260 45.570 ;
        RECT 110.680 80.350 115.130 80.770 ;
        RECT 110.680 44.110 111.100 80.350 ;
        RECT 114.900 79.700 115.130 80.350 ;
        RECT 115.390 81.740 115.620 84.700 ;
        RECT 115.390 80.460 118.660 81.740 ;
        RECT 115.390 79.700 115.620 80.460 ;
        RECT 103.250 43.690 111.100 44.110 ;
        RECT 103.250 38.590 103.670 43.690 ;
        RECT 81.810 37.870 106.840 38.590 ;
        RECT 105.920 37.625 106.840 37.870 ;
        RECT 105.885 36.730 106.880 37.625 ;
        RECT 58.920 35.300 59.380 35.660 ;
        RECT 58.920 31.970 59.380 32.330 ;
        RECT 58.970 31.660 59.330 31.970 ;
        RECT 60.780 31.660 61.010 33.380 ;
        RECT 58.970 31.300 61.010 31.660 ;
        RECT 60.780 29.380 61.010 31.300 ;
        RECT 105.870 29.095 106.880 30.005 ;
        RECT 105.920 27.070 106.830 29.095 ;
        RECT 110.660 27.070 110.890 33.380 ;
        RECT 105.920 26.160 110.890 27.070 ;
        RECT 110.660 17.380 110.890 26.160 ;
      LAYER via ;
        RECT 65.940 69.660 66.480 70.200 ;
        RECT 81.790 69.615 82.740 70.565 ;
        RECT 195.705 109.110 196.115 109.520 ;
        RECT 202.120 109.120 202.520 109.520 ;
        RECT 65.950 63.860 66.490 64.400 ;
        RECT 81.810 61.770 82.730 62.690 ;
        RECT 79.815 56.560 80.185 56.930 ;
        RECT 44.850 45.290 45.110 45.550 ;
        RECT 48.880 45.290 49.140 45.550 ;
        RECT 57.060 45.290 57.320 45.550 ;
        RECT 60.265 45.265 60.570 45.570 ;
        RECT 77.365 45.260 77.675 45.570 ;
        RECT 85.320 56.580 85.665 56.925 ;
        RECT 84.030 45.250 84.350 45.570 ;
        RECT 117.330 80.460 118.610 81.740 ;
        RECT 105.935 36.730 106.830 37.625 ;
        RECT 58.970 35.300 59.330 35.660 ;
        RECT 58.970 31.970 59.330 32.330 ;
        RECT 105.920 29.095 106.830 30.005 ;
      LAYER met2 ;
        RECT 195.705 109.520 196.115 109.570 ;
        RECT 202.120 109.520 202.520 109.570 ;
        RECT 195.705 109.110 202.520 109.520 ;
        RECT 195.705 109.060 196.115 109.110 ;
        RECT 202.120 109.070 202.520 109.110 ;
        RECT 117.330 81.780 118.610 81.790 ;
        RECT 119.320 81.780 120.660 81.820 ;
        RECT 117.310 80.440 120.660 81.780 ;
        RECT 117.330 80.430 120.660 80.440 ;
        RECT 117.330 80.410 118.610 80.430 ;
        RECT 119.320 80.380 120.660 80.430 ;
        RECT 65.940 64.450 66.480 70.250 ;
        RECT 65.940 63.850 66.490 64.450 ;
        RECT 65.950 63.810 66.490 63.850 ;
        RECT 81.790 61.730 82.740 70.615 ;
        RECT 81.810 61.720 82.730 61.730 ;
        RECT 79.815 56.930 80.185 56.980 ;
        RECT 85.320 56.930 85.665 56.975 ;
        RECT 79.815 56.560 85.670 56.930 ;
        RECT 79.815 56.510 80.185 56.560 ;
        RECT 85.320 56.530 85.665 56.560 ;
        RECT 44.850 45.550 45.110 45.600 ;
        RECT 48.880 45.550 49.140 45.600 ;
        RECT 44.850 45.290 49.140 45.550 ;
        RECT 44.850 45.240 45.110 45.290 ;
        RECT 48.880 45.240 49.140 45.290 ;
        RECT 57.060 45.570 57.320 45.600 ;
        RECT 60.265 45.570 60.570 45.620 ;
        RECT 77.365 45.570 77.675 45.620 ;
        RECT 84.030 45.570 84.350 45.620 ;
        RECT 57.060 45.265 60.570 45.570 ;
        RECT 57.060 45.240 57.320 45.265 ;
        RECT 60.265 45.215 60.570 45.265 ;
        RECT 77.360 45.250 84.350 45.570 ;
        RECT 77.365 45.210 77.675 45.250 ;
        RECT 84.030 45.200 84.350 45.250 ;
        RECT 58.970 31.920 59.330 35.710 ;
        RECT 105.935 30.900 106.830 37.675 ;
        RECT 105.920 29.045 106.830 30.900 ;
      LAYER via2 ;
        RECT 119.320 80.430 120.660 81.770 ;
      LAYER met3 ;
        RECT 119.290 81.795 121.390 81.810 ;
        RECT 119.270 81.790 121.390 81.795 ;
        RECT 119.270 80.405 122.750 81.790 ;
        RECT 119.290 80.380 122.750 80.405 ;
      LAYER via3 ;
        RECT 121.290 80.380 122.700 81.790 ;
      LAYER met4 ;
        RECT 132.625 85.735 156.895 115.345 ;
        RECT 160.625 85.735 184.895 115.345 ;
        RECT 141.140 83.200 148.240 85.735 ;
        RECT 169.140 83.200 176.240 85.735 ;
        RECT 141.140 81.860 176.240 83.200 ;
        RECT 122.700 81.820 176.240 81.860 ;
        RECT 121.270 80.380 176.240 81.820 ;
        RECT 121.285 80.375 122.705 80.380 ;
        RECT 141.140 79.060 176.240 80.380 ;
        RECT 141.140 77.345 148.240 79.060 ;
        RECT 169.140 77.345 176.240 79.060 ;
        RECT 132.625 47.735 156.895 77.345 ;
        RECT 160.625 47.735 184.895 77.345 ;
  END
END tt_um_keremergunay_two_stage_opamp
END LIBRARY


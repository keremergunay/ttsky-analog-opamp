VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_keremergunay_two_stage_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_keremergunay_two_stage_opamp ;
  ORIGIN 0.000 0.010 ;
  SIZE 219.600 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 142.830 224.750 143.130 225.750 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 145.590 224.750 145.890 225.750 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.070 224.750 140.370 225.750 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER li1 ;
        RECT 72.580 63.010 73.580 63.180 ;
      LAYER mcon ;
        RECT 72.660 63.010 73.500 63.180 ;
      LAYER met1 ;
        RECT 71.550 65.400 74.260 65.450 ;
        RECT 71.550 64.460 74.710 65.400 ;
        RECT 71.550 64.420 74.260 64.460 ;
        RECT 72.550 63.950 73.550 64.420 ;
        RECT 72.930 63.210 73.250 63.950 ;
        RECT 72.600 62.980 73.560 63.210 ;
      LAYER via ;
        RECT 73.720 64.460 74.660 65.400 ;
      LAYER met2 ;
        RECT 73.720 65.410 74.660 65.450 ;
        RECT 75.040 65.410 75.960 65.420 ;
        RECT 73.720 64.450 75.970 65.410 ;
        RECT 73.720 64.410 74.660 64.450 ;
        RECT 75.040 64.400 75.960 64.450 ;
      LAYER via2 ;
        RECT 75.040 64.450 75.960 65.370 ;
      LAYER met3 ;
        RECT 74.990 65.370 76.010 65.395 ;
        RECT 74.990 64.470 77.470 65.370 ;
        RECT 74.990 64.450 77.420 64.470 ;
        RECT 74.990 64.425 76.010 64.450 ;
      LAYER via3 ;
        RECT 76.520 64.470 77.420 65.370 ;
      LAYER met4 ;
        RECT 76.515 65.370 77.425 65.375 ;
        RECT 76.515 64.470 125.230 65.370 ;
        RECT 76.515 64.465 77.425 64.470 ;
        RECT 124.330 43.390 125.230 64.470 ;
        RECT 124.330 42.490 151.710 43.390 ;
        RECT 150.810 -0.010 151.710 42.490 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER li1 ;
        RECT 50.790 62.970 51.790 63.140 ;
      LAYER mcon ;
        RECT 50.870 62.970 51.710 63.140 ;
      LAYER met1 ;
        RECT 49.780 65.020 53.260 65.030 ;
        RECT 49.780 64.970 54.120 65.020 ;
        RECT 49.780 64.030 54.570 64.970 ;
        RECT 50.770 64.010 51.770 64.030 ;
        RECT 51.150 63.170 51.430 64.010 ;
        RECT 52.900 63.990 54.120 64.030 ;
        RECT 50.810 62.940 51.770 63.170 ;
      LAYER via ;
        RECT 53.580 64.030 54.520 64.970 ;
      LAYER met2 ;
        RECT 53.580 64.980 54.520 65.020 ;
        RECT 54.900 64.980 55.820 64.990 ;
        RECT 53.580 64.020 55.830 64.980 ;
        RECT 53.580 63.980 54.520 64.020 ;
        RECT 54.900 63.970 55.820 64.020 ;
      LAYER via2 ;
        RECT 54.900 64.020 55.820 64.940 ;
      LAYER met3 ;
        RECT 54.850 64.940 55.870 64.965 ;
        RECT 54.850 64.040 57.330 64.940 ;
        RECT 54.850 64.020 57.280 64.040 ;
        RECT 54.850 63.995 55.870 64.020 ;
      LAYER via3 ;
        RECT 56.380 64.040 57.280 64.940 ;
      LAYER met4 ;
        RECT 57.230 64.945 62.880 64.990 ;
        RECT 56.375 64.090 62.880 64.945 ;
        RECT 56.375 64.040 57.850 64.090 ;
        RECT 56.375 64.035 57.285 64.040 ;
        RECT 61.980 55.290 62.880 64.090 ;
        RECT 61.980 54.390 118.690 55.290 ;
        RECT 117.790 39.540 118.690 54.390 ;
        RECT 117.790 38.640 132.390 39.540 ;
        RECT 131.490 -0.010 132.390 38.640 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 11.710199 ;
    PORT
      LAYER li1 ;
        RECT 209.430 110.770 209.600 135.190 ;
        RECT 207.080 17.370 207.250 33.410 ;
      LAYER mcon ;
        RECT 209.430 110.850 209.600 135.110 ;
        RECT 207.080 17.450 207.250 33.330 ;
      LAYER met1 ;
        RECT 209.400 120.385 209.630 135.170 ;
        RECT 197.305 118.535 209.630 120.385 ;
        RECT 197.305 83.520 199.155 118.535 ;
        RECT 209.400 110.790 209.630 118.535 ;
        RECT 217.330 90.245 218.440 90.250 ;
        RECT 217.320 89.255 218.440 90.245 ;
        RECT 197.305 83.090 203.360 83.520 ;
        RECT 192.470 82.540 203.360 83.090 ;
        RECT 192.470 81.240 199.155 82.540 ;
        RECT 202.380 82.210 203.360 82.540 ;
        RECT 217.330 82.210 218.440 89.255 ;
        RECT 218.600 82.210 219.600 82.250 ;
        RECT 202.380 81.250 219.600 82.210 ;
        RECT 192.530 81.190 194.530 81.240 ;
        RECT 202.380 81.230 219.030 81.250 ;
        RECT 202.380 35.580 203.360 81.230 ;
        RECT 202.330 34.620 203.390 35.580 ;
        RECT 202.380 34.610 203.360 34.620 ;
        RECT 202.335 28.905 203.365 29.835 ;
        RECT 202.385 25.500 203.315 28.905 ;
        RECT 207.050 25.500 207.280 33.390 ;
        RECT 202.385 24.570 207.280 25.500 ;
        RECT 207.050 17.390 207.280 24.570 ;
      LAYER via ;
        RECT 217.370 89.255 218.360 90.245 ;
        RECT 192.580 81.190 194.480 83.090 ;
        RECT 202.380 34.620 203.340 35.580 ;
        RECT 202.385 28.905 203.315 29.835 ;
      LAYER met2 ;
        RECT 217.410 91.940 218.350 91.980 ;
        RECT 217.370 89.205 218.360 91.940 ;
        RECT 189.100 83.090 190.950 83.140 ;
        RECT 192.580 83.090 194.480 83.140 ;
        RECT 189.050 81.190 194.480 83.090 ;
        RECT 192.580 81.140 194.480 81.190 ;
        RECT 202.380 29.840 203.340 35.630 ;
        RECT 202.380 28.890 203.330 29.840 ;
        RECT 202.385 28.855 203.315 28.890 ;
      LAYER via2 ;
        RECT 217.410 90.990 218.350 91.930 ;
        RECT 189.100 81.240 190.950 83.090 ;
      LAYER met3 ;
        RECT 131.690 116.020 185.940 116.190 ;
        RECT 131.690 115.590 186.075 116.020 ;
        RECT 131.690 85.300 158.075 115.590 ;
        RECT 131.860 85.020 158.075 85.300 ;
        RECT 159.920 85.020 186.075 115.590 ;
        RECT 217.410 93.510 218.350 93.520 ;
        RECT 217.370 92.610 218.370 93.510 ;
        RECT 217.410 91.955 218.350 92.610 ;
        RECT 217.360 90.965 218.400 91.955 ;
        RECT 131.860 78.020 132.460 85.020 ;
        RECT 185.340 83.090 185.940 85.020 ;
        RECT 189.050 83.090 191.000 83.115 ;
        RECT 185.290 81.240 191.000 83.090 ;
        RECT 185.340 78.020 185.940 81.240 ;
        RECT 189.050 81.215 191.000 81.240 ;
        RECT 131.860 47.450 158.075 78.020 ;
        RECT 159.920 47.450 186.075 78.020 ;
        RECT 131.860 47.020 186.075 47.450 ;
        RECT 131.860 46.850 186.060 47.020 ;
      LAYER via3 ;
        RECT 157.655 85.160 157.975 115.880 ;
        RECT 185.655 85.160 185.975 115.880 ;
        RECT 217.420 92.610 218.320 93.510 ;
        RECT 157.655 47.160 157.975 77.880 ;
        RECT 185.655 47.160 185.975 77.880 ;
      LAYER met4 ;
        RECT 33.000 134.960 202.140 135.860 ;
        RECT 33.000 42.600 33.900 134.960 ;
        RECT 157.575 85.080 158.055 115.960 ;
        RECT 185.575 85.080 186.055 115.960 ;
        RECT 201.240 115.260 202.140 134.960 ;
        RECT 201.240 114.360 204.220 115.260 ;
        RECT 203.320 93.510 204.220 114.360 ;
        RECT 217.415 93.510 218.325 93.515 ;
        RECT 203.320 92.610 218.325 93.510 ;
        RECT 217.415 92.605 218.325 92.610 ;
        RECT 157.575 47.080 158.055 77.960 ;
        RECT 185.575 47.080 186.055 77.960 ;
        RECT 33.000 41.700 87.120 42.600 ;
        RECT 86.220 12.750 87.120 41.700 ;
        RECT 86.220 11.850 113.070 12.750 ;
        RECT 112.170 -0.010 113.070 11.850 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 29.000000 ;
    ANTENNADIFFAREA 1.740000 ;
    PORT
      LAYER li1 ;
        RECT 26.435 41.370 26.605 41.870 ;
        RECT 24.180 41.140 26.220 41.310 ;
        RECT 18.015 33.525 18.515 33.695 ;
        RECT 32.225 33.455 32.725 33.625 ;
        RECT 61.030 33.550 61.530 33.720 ;
        RECT 110.910 33.550 111.410 33.720 ;
        RECT 207.310 33.580 208.310 33.750 ;
        RECT 17.785 31.315 17.955 33.355 ;
        RECT 31.995 31.245 32.165 33.285 ;
      LAYER mcon ;
        RECT 26.435 41.450 26.605 41.790 ;
        RECT 24.260 41.140 26.140 41.310 ;
        RECT 18.095 33.525 18.435 33.695 ;
        RECT 32.305 33.455 32.645 33.625 ;
        RECT 61.110 33.550 61.450 33.720 ;
        RECT 110.990 33.550 111.330 33.720 ;
        RECT 207.390 33.580 208.230 33.750 ;
        RECT 17.785 31.395 17.955 33.275 ;
        RECT 31.995 31.325 32.165 33.205 ;
      LAYER met1 ;
        RECT 26.405 41.760 26.635 41.850 ;
        RECT 26.405 41.390 26.710 41.760 ;
        RECT 24.200 41.110 26.200 41.340 ;
        RECT 24.940 39.790 25.180 41.110 ;
        RECT 26.470 39.790 26.710 41.390 ;
        RECT 24.940 39.550 26.710 39.790 ;
        RECT 13.250 34.290 14.270 34.410 ;
        RECT 14.790 34.290 15.790 34.360 ;
        RECT 13.250 33.780 15.790 34.290 ;
        RECT 24.940 33.780 25.180 39.550 ;
        RECT 13.250 33.550 208.290 33.780 ;
        RECT 13.250 33.540 208.260 33.550 ;
        RECT 13.250 33.360 15.790 33.540 ;
        RECT 13.250 33.270 15.370 33.360 ;
        RECT 13.250 24.475 14.270 33.270 ;
        RECT 16.620 32.520 16.890 33.540 ;
        RECT 18.035 33.495 18.495 33.540 ;
        RECT 17.755 32.520 17.985 33.335 ;
        RECT 16.620 32.250 17.985 32.520 ;
        RECT 30.460 32.620 30.700 33.540 ;
        RECT 32.245 33.425 32.705 33.540 ;
        RECT 61.050 33.520 61.510 33.540 ;
        RECT 110.930 33.520 111.390 33.540 ;
        RECT 31.965 32.620 32.195 33.265 ;
        RECT 30.460 32.380 32.195 32.620 ;
        RECT 17.755 31.335 17.985 32.250 ;
        RECT 31.965 31.265 32.195 32.380 ;
        RECT 13.240 23.545 14.270 24.475 ;
        RECT 13.250 23.540 14.270 23.545 ;
      LAYER via ;
        RECT 13.290 23.545 14.220 24.475 ;
      LAYER met2 ;
        RECT 13.290 23.660 14.220 24.525 ;
        RECT 13.270 22.780 14.220 23.660 ;
        RECT 13.270 21.780 14.230 22.780 ;
        RECT 13.290 21.740 14.230 21.780 ;
      LAYER via2 ;
        RECT 13.290 21.790 14.230 22.730 ;
      LAYER met3 ;
        RECT 13.240 21.765 14.280 22.755 ;
        RECT 13.290 21.170 14.230 21.765 ;
        RECT 13.220 20.270 14.230 21.170 ;
        RECT 13.290 20.230 14.230 20.270 ;
      LAYER via3 ;
        RECT 13.270 20.270 14.170 21.170 ;
      LAYER met4 ;
        RECT 13.265 20.265 14.175 21.175 ;
        RECT 13.270 19.950 14.170 20.265 ;
        RECT 13.270 19.050 82.830 19.950 ;
        RECT 81.930 3.330 82.830 19.050 ;
        RECT 81.930 2.430 93.750 3.330 ;
        RECT 92.850 -0.010 93.750 2.430 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.530 -0.010 74.430 0.990 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.210 -0.010 55.110 0.990 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.890 -0.010 35.790 0.990 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.570 -0.010 16.470 0.990 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 137.310 224.750 137.610 225.750 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.550 224.750 134.850 225.750 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 131.790 224.750 132.090 225.750 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.030 224.750 129.330 225.750 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 126.270 224.750 126.570 225.750 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 123.510 224.750 123.810 225.750 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 120.750 224.750 121.050 225.750 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.990 224.750 118.290 225.750 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 115.230 224.750 115.530 225.750 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.470 224.750 112.770 225.750 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 109.710 224.750 110.010 225.750 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.950 224.750 107.250 225.750 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 104.190 224.750 104.490 225.750 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 101.430 224.750 101.730 225.750 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.670 224.750 98.970 225.750 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.910 224.750 96.210 225.750 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.990 224.750 49.290 225.750 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.230 224.750 46.530 225.750 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 43.470 224.750 43.770 225.750 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.710 224.750 41.010 225.750 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.950 224.750 38.250 225.750 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.190 224.750 35.490 225.750 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.430 224.750 32.730 225.750 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.670 224.750 29.970 225.750 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 71.070 224.750 71.370 225.750 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.310 224.750 68.610 225.750 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 65.550 224.750 65.850 225.750 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.790 224.750 63.090 225.750 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 60.030 224.750 60.330 225.750 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 57.270 224.750 57.570 225.750 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.510 224.750 54.810 225.750 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.750 224.750 52.050 225.750 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.150 224.750 93.450 225.750 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.390 224.750 90.690 225.750 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 87.630 224.750 87.930 225.750 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.870 224.750 85.170 225.750 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 82.110 224.750 82.410 225.750 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 79.350 224.750 79.650 225.750 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 76.590 224.750 76.890 225.750 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.830 224.750 74.130 225.750 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 47.890 70.460 54.850 132.300 ;
        RECT 69.470 70.430 76.430 132.270 ;
        RECT 89.960 111.330 92.420 118.170 ;
        RECT 208.680 109.690 211.140 135.910 ;
        RECT 23.460 53.100 27.300 55.560 ;
        RECT 23.390 46.970 27.230 49.430 ;
        RECT 23.460 40.390 27.300 42.850 ;
      LAYER li1 ;
        RECT 209.260 135.560 210.560 135.730 ;
        RECT 48.470 131.950 54.270 132.120 ;
        RECT 70.050 131.920 75.850 132.090 ;
        RECT 53.930 71.540 54.100 131.580 ;
        RECT 75.510 71.510 75.680 131.550 ;
        RECT 90.540 117.820 91.840 117.990 ;
        RECT 91.500 112.410 91.670 117.450 ;
        RECT 210.220 110.770 210.390 135.190 ;
        RECT 23.640 53.680 23.810 54.980 ;
        RECT 24.180 54.640 26.220 54.810 ;
        RECT 23.570 47.550 23.740 48.850 ;
        RECT 23.640 40.970 23.810 42.270 ;
      LAYER mcon ;
        RECT 209.340 135.560 210.480 135.730 ;
        RECT 48.550 131.950 54.190 132.120 ;
        RECT 70.130 131.920 75.770 132.090 ;
        RECT 53.930 71.620 54.100 131.500 ;
        RECT 75.510 71.590 75.680 131.470 ;
        RECT 90.620 117.820 91.760 117.990 ;
        RECT 91.500 112.490 91.670 117.370 ;
        RECT 210.220 110.850 210.390 135.110 ;
        RECT 23.640 53.760 23.810 54.900 ;
        RECT 24.260 54.640 26.140 54.810 ;
        RECT 23.570 47.630 23.740 48.770 ;
        RECT 23.640 41.050 23.810 42.190 ;
      LAYER met1 ;
        RECT 60.200 161.860 62.270 161.865 ;
        RECT 60.170 159.895 62.270 161.860 ;
        RECT 60.170 142.780 62.250 159.895 ;
        RECT 60.225 138.385 62.200 142.780 ;
        RECT 22.540 138.095 212.465 138.385 ;
        RECT 22.540 56.765 22.830 138.095 ;
        RECT 50.955 132.150 51.245 138.095 ;
        RECT 48.490 131.920 54.250 132.150 ;
        RECT 53.900 119.335 54.130 131.560 ;
        RECT 57.145 119.335 57.435 138.095 ;
        RECT 61.080 137.470 62.080 138.095 ;
        RECT 72.815 135.275 73.105 138.095 ;
        RECT 72.815 134.985 79.505 135.275 ;
        RECT 72.815 132.120 73.105 134.985 ;
        RECT 70.070 131.890 75.830 132.120 ;
        RECT 53.900 119.045 57.435 119.335 ;
        RECT 75.480 126.365 75.710 131.530 ;
        RECT 79.215 126.365 79.505 134.985 ;
        RECT 75.480 126.075 79.505 126.365 ;
        RECT 53.900 71.560 54.130 119.045 ;
        RECT 75.480 71.530 75.710 126.075 ;
        RECT 90.955 118.905 91.245 138.095 ;
        RECT 209.675 135.760 209.965 138.095 ;
        RECT 209.280 135.530 210.540 135.760 ;
        RECT 210.190 129.785 210.420 135.170 ;
        RECT 212.175 129.785 212.465 138.095 ;
        RECT 210.190 129.495 212.465 129.785 ;
        RECT 90.955 118.615 94.045 118.905 ;
        RECT 90.955 118.020 91.245 118.615 ;
        RECT 90.560 117.790 91.820 118.020 ;
        RECT 91.470 115.155 91.700 117.430 ;
        RECT 93.755 115.155 94.045 118.615 ;
        RECT 91.470 114.865 94.045 115.155 ;
        RECT 91.470 112.430 91.700 114.865 ;
        RECT 210.190 110.790 210.420 129.495 ;
        RECT 22.540 56.475 25.155 56.765 ;
        RECT 22.540 54.465 22.830 56.475 ;
        RECT 23.610 54.465 23.840 54.960 ;
        RECT 24.865 54.840 25.155 56.475 ;
        RECT 24.200 54.610 26.200 54.840 ;
        RECT 22.540 54.175 23.840 54.465 ;
        RECT 22.540 48.385 22.830 54.175 ;
        RECT 23.610 53.700 23.840 54.175 ;
        RECT 23.540 48.385 23.770 48.830 ;
        RECT 22.540 48.095 23.770 48.385 ;
        RECT 22.540 41.690 22.830 48.095 ;
        RECT 23.540 47.570 23.770 48.095 ;
        RECT 23.610 41.690 23.840 42.250 ;
        RECT 22.540 41.400 23.840 41.690 ;
        RECT 23.610 40.990 23.840 41.400 ;
      LAYER via ;
        RECT 60.250 159.895 62.220 161.865 ;
      LAYER met2 ;
        RECT 60.250 162.990 62.230 165.050 ;
        RECT 60.250 159.845 62.220 162.990 ;
      LAYER via2 ;
        RECT 60.270 163.040 62.230 165.000 ;
      LAYER met3 ;
        RECT 60.270 168.690 62.230 168.730 ;
        RECT 60.230 166.690 62.330 168.690 ;
        RECT 60.270 165.025 62.230 166.690 ;
        RECT 60.220 163.015 62.280 165.025 ;
      LAYER via3 ;
        RECT 60.280 166.690 62.280 168.690 ;
      LAYER met4 ;
        RECT 0.000 221.910 22.930 223.910 ;
        RECT 0.000 4.990 2.000 221.910 ;
        RECT 20.930 172.960 22.930 221.910 ;
        RECT 20.930 170.960 62.280 172.960 ;
        RECT 60.280 168.695 62.280 170.960 ;
        RECT 60.275 166.685 62.285 168.695 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 114.170 78.940 116.330 85.730 ;
        RECT 49.810 59.040 52.770 63.830 ;
        RECT 71.600 59.080 74.560 63.870 ;
        RECT 17.035 30.595 19.495 34.385 ;
        RECT 31.245 30.525 33.705 34.315 ;
        RECT 60.050 28.620 62.510 34.410 ;
        RECT 109.930 16.620 112.390 34.410 ;
        RECT 206.330 16.650 209.290 34.440 ;
      LAYER li1 ;
        RECT 114.750 79.120 115.750 79.290 ;
        RECT 50.390 59.220 52.190 59.390 ;
        RECT 72.180 59.260 73.980 59.430 ;
        RECT 18.575 31.315 18.745 33.355 ;
        RECT 32.785 31.245 32.955 33.285 ;
        RECT 17.615 30.775 18.915 30.945 ;
        RECT 31.825 30.705 33.125 30.875 ;
        RECT 61.590 29.340 61.760 33.380 ;
        RECT 60.630 28.800 61.930 28.970 ;
        RECT 111.470 17.340 111.640 33.380 ;
        RECT 208.370 17.370 208.540 33.410 ;
        RECT 110.510 16.800 111.810 16.970 ;
        RECT 206.910 16.830 208.710 17.000 ;
      LAYER mcon ;
        RECT 114.830 79.120 115.670 79.290 ;
        RECT 50.470 59.220 52.110 59.390 ;
        RECT 72.260 59.260 73.900 59.430 ;
        RECT 18.575 31.395 18.745 33.275 ;
        RECT 32.785 31.325 32.955 33.205 ;
        RECT 17.695 30.775 18.835 30.945 ;
        RECT 31.905 30.705 33.045 30.875 ;
        RECT 61.590 29.420 61.760 33.300 ;
        RECT 60.710 28.800 61.850 28.970 ;
        RECT 111.470 17.420 111.640 33.300 ;
        RECT 208.370 17.450 208.540 33.330 ;
        RECT 110.590 16.800 111.730 16.970 ;
        RECT 206.990 16.830 208.630 17.000 ;
      LAYER met1 ;
        RECT 114.770 79.090 115.730 79.320 ;
        RECT 50.410 59.190 52.170 59.420 ;
        RECT 72.200 59.230 73.960 59.460 ;
        RECT 51.280 55.360 51.640 59.190 ;
        RECT 72.955 58.320 73.345 59.230 ;
        RECT 72.955 57.930 73.840 58.320 ;
        RECT 73.450 57.215 73.840 57.930 ;
        RECT 73.425 56.860 73.880 57.215 ;
        RECT 73.450 56.850 73.840 56.860 ;
        RECT 47.580 55.000 51.640 55.360 ;
        RECT 47.580 34.480 47.940 55.000 ;
        RECT 115.070 37.115 115.420 79.090 ;
        RECT 115.070 36.765 144.845 37.115 ;
        RECT 144.495 35.605 144.845 36.765 ;
        RECT 144.445 35.255 144.895 35.605 ;
        RECT 47.530 34.120 47.990 34.480 ;
        RECT 18.545 31.800 18.775 33.335 ;
        RECT 32.755 32.120 32.985 33.265 ;
        RECT 18.545 31.335 18.800 31.800 ;
        RECT 18.590 30.975 18.800 31.335 ;
        RECT 32.755 31.760 36.270 32.120 ;
        RECT 32.755 31.265 32.985 31.760 ;
        RECT 17.635 30.745 18.895 30.975 ;
        RECT 18.170 10.200 18.530 30.745 ;
        RECT 31.845 30.675 33.105 30.905 ;
        RECT 31.980 10.200 32.340 30.675 ;
        RECT 35.910 10.200 36.270 31.760 ;
        RECT 47.530 31.720 47.990 32.080 ;
        RECT 47.580 10.200 47.940 31.720 ;
        RECT 61.560 31.640 61.790 33.360 ;
        RECT 73.420 31.830 73.880 32.190 ;
        RECT 61.560 31.280 64.140 31.640 ;
        RECT 61.560 29.360 61.790 31.280 ;
        RECT 60.650 28.770 61.910 29.000 ;
        RECT 60.940 27.610 61.300 28.770 ;
        RECT 63.780 27.610 64.140 31.280 ;
        RECT 60.940 27.250 64.140 27.610 ;
        RECT 60.940 10.200 61.300 27.250 ;
        RECT 73.470 10.200 73.830 31.830 ;
        RECT 111.440 27.610 111.670 33.360 ;
        RECT 144.490 33.160 144.850 33.170 ;
        RECT 144.440 32.800 144.900 33.160 ;
        RECT 111.440 27.250 114.450 27.610 ;
        RECT 111.440 17.360 111.670 27.250 ;
        RECT 110.530 16.770 111.790 17.000 ;
        RECT 110.850 15.840 111.210 16.770 ;
        RECT 114.090 15.840 114.450 27.250 ;
        RECT 110.850 15.480 114.450 15.840 ;
        RECT 75.380 10.470 76.380 10.530 ;
        RECT 74.370 10.200 76.380 10.470 ;
        RECT 110.850 10.200 111.210 15.480 ;
        RECT 144.490 10.200 144.850 32.800 ;
        RECT 208.340 25.130 208.570 33.390 ;
        RECT 208.340 24.770 211.810 25.130 ;
        RECT 208.340 17.390 208.570 24.770 ;
        RECT 206.930 16.800 208.690 17.030 ;
        RECT 207.400 15.010 207.760 16.800 ;
        RECT 211.450 15.010 211.810 24.770 ;
        RECT 207.400 14.650 211.810 15.010 ;
        RECT 207.400 10.200 207.760 14.650 ;
        RECT 18.170 9.840 207.760 10.200 ;
        RECT 74.370 9.530 76.380 9.840 ;
        RECT 74.370 8.630 75.435 9.530 ;
        RECT 74.370 7.565 76.495 8.630 ;
        RECT 75.430 7.180 76.495 7.565 ;
        RECT 72.630 4.940 77.080 7.180 ;
      LAYER via ;
        RECT 73.475 56.860 73.830 57.215 ;
        RECT 144.495 35.255 144.845 35.605 ;
        RECT 47.580 34.120 47.940 34.480 ;
        RECT 47.580 31.720 47.940 32.080 ;
        RECT 73.470 31.830 73.830 32.190 ;
        RECT 144.490 32.800 144.850 33.160 ;
        RECT 72.710 5.025 74.805 7.120 ;
      LAYER met2 ;
        RECT 47.580 31.670 47.940 34.530 ;
        RECT 73.475 32.530 73.830 57.265 ;
        RECT 144.495 35.620 144.845 35.655 ;
        RECT 144.490 32.750 144.850 35.620 ;
        RECT 73.470 31.830 73.840 32.530 ;
        RECT 73.470 31.780 73.830 31.830 ;
        RECT 72.710 7.120 74.805 7.170 ;
        RECT 70.625 7.080 74.805 7.120 ;
        RECT 68.600 5.030 74.805 7.080 ;
        RECT 68.600 4.940 70.750 5.030 ;
        RECT 72.680 5.025 74.805 5.030 ;
        RECT 72.710 4.975 74.805 5.025 ;
        RECT 68.600 4.900 70.680 4.940 ;
      LAYER via2 ;
        RECT 68.600 4.950 70.680 7.030 ;
      LAYER met3 ;
        RECT 68.550 7.030 70.730 7.055 ;
        RECT 65.100 4.925 70.730 7.030 ;
        RECT 65.100 4.880 69.280 4.925 ;
      LAYER via3 ;
        RECT 65.200 4.990 67.200 6.990 ;
      LAYER met4 ;
        RECT 3.000 6.990 5.000 220.750 ;
        RECT 65.195 6.990 67.205 6.995 ;
        RECT 3.000 4.990 67.205 6.990 ;
        RECT 65.195 4.985 67.205 4.990 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 48.640 71.540 48.810 131.580 ;
        RECT 70.220 71.510 70.390 131.550 ;
        RECT 90.710 112.410 90.880 117.450 ;
        RECT 90.940 112.025 91.440 112.195 ;
        RECT 209.660 110.385 210.160 110.555 ;
        RECT 115.085 84.870 115.415 85.040 ;
        RECT 114.920 79.660 115.090 84.700 ;
        RECT 115.410 79.660 115.580 84.700 ;
        RECT 48.870 71.155 53.870 71.325 ;
        RECT 70.450 71.125 75.450 71.295 ;
        RECT 50.560 59.760 50.730 62.800 ;
        RECT 51.850 59.760 52.020 62.800 ;
        RECT 72.350 59.800 72.520 62.840 ;
        RECT 73.640 59.800 73.810 62.840 ;
        RECT 26.435 54.080 26.605 54.580 ;
        RECT 24.180 53.850 26.220 54.020 ;
        RECT 24.110 48.510 26.150 48.680 ;
        RECT 26.365 47.950 26.535 48.450 ;
        RECT 24.110 47.720 26.150 47.890 ;
        RECT 24.180 41.930 26.220 42.100 ;
        RECT 60.800 29.340 60.970 33.380 ;
        RECT 110.680 17.340 110.850 33.380 ;
      LAYER mcon ;
        RECT 48.640 71.620 48.810 131.500 ;
        RECT 70.220 71.590 70.390 131.470 ;
        RECT 90.710 112.490 90.880 117.370 ;
        RECT 91.020 112.025 91.360 112.195 ;
        RECT 209.740 110.385 210.080 110.555 ;
        RECT 115.165 84.870 115.335 85.040 ;
        RECT 114.920 79.740 115.090 84.620 ;
        RECT 115.410 79.740 115.580 84.620 ;
        RECT 48.950 71.155 53.790 71.325 ;
        RECT 70.530 71.125 75.370 71.295 ;
        RECT 50.560 59.840 50.730 62.720 ;
        RECT 51.850 59.840 52.020 62.720 ;
        RECT 72.350 59.880 72.520 62.760 ;
        RECT 73.640 59.880 73.810 62.760 ;
        RECT 26.435 54.160 26.605 54.500 ;
        RECT 24.260 53.850 26.140 54.020 ;
        RECT 24.190 48.510 26.070 48.680 ;
        RECT 26.365 48.030 26.535 48.370 ;
        RECT 24.190 47.720 26.070 47.890 ;
        RECT 24.260 41.930 26.140 42.100 ;
        RECT 60.800 29.420 60.970 33.300 ;
        RECT 110.680 17.420 110.850 33.300 ;
      LAYER met1 ;
        RECT 48.610 82.700 48.840 131.560 ;
        RECT 43.140 82.200 48.840 82.700 ;
        RECT 43.140 68.170 43.640 82.200 ;
        RECT 48.610 71.560 48.840 82.200 ;
        RECT 70.190 74.245 70.420 131.530 ;
        RECT 101.250 120.835 190.865 121.180 ;
        RECT 90.680 114.580 90.910 117.430 ;
        RECT 65.920 73.675 70.420 74.245 ;
        RECT 48.890 71.125 53.850 71.355 ;
        RECT 50.950 68.170 51.450 71.125 ;
        RECT 65.920 70.180 66.490 73.675 ;
        RECT 70.190 71.530 70.420 73.675 ;
        RECT 81.770 113.620 90.910 114.580 ;
        RECT 70.470 71.095 75.430 71.325 ;
        RECT 65.880 69.640 66.520 70.180 ;
        RECT 72.770 68.170 73.270 71.095 ;
        RECT 81.770 70.545 82.730 113.620 ;
        RECT 90.680 112.430 90.910 113.620 ;
        RECT 90.960 112.170 91.420 112.225 ;
        RECT 90.960 111.995 91.470 112.170 ;
        RECT 90.970 103.150 91.470 111.995 ;
        RECT 85.860 102.650 91.470 103.150 ;
        RECT 81.730 69.595 82.780 70.545 ;
        RECT 81.770 69.580 82.730 69.595 ;
        RECT 85.860 68.170 86.360 102.650 ;
        RECT 101.250 95.215 101.595 120.835 ;
        RECT 190.520 109.470 190.865 120.835 ;
        RECT 209.680 110.355 210.140 110.585 ;
        RECT 209.720 109.500 210.120 110.355 ;
        RECT 195.350 109.470 196.155 109.500 ;
        RECT 190.520 109.125 196.155 109.470 ;
        RECT 195.350 109.090 196.155 109.125 ;
        RECT 202.060 109.100 210.120 109.500 ;
        RECT 195.350 109.080 196.110 109.090 ;
        RECT 43.140 67.670 86.360 68.170 ;
        RECT 90.720 94.870 101.595 95.215 ;
        RECT 43.140 61.280 43.640 67.670 ;
        RECT 69.695 66.015 79.590 66.405 ;
        RECT 65.890 63.840 66.530 64.380 ;
        RECT 50.530 61.280 50.760 62.780 ;
        RECT 43.140 60.780 50.760 61.280 ;
        RECT 50.530 59.780 50.760 60.780 ;
        RECT 51.820 61.250 52.050 62.780 ;
        RECT 65.940 61.420 66.480 63.840 ;
        RECT 69.695 61.420 70.085 66.015 ;
        RECT 72.320 61.420 72.550 62.820 ;
        RECT 51.820 60.890 59.320 61.250 ;
        RECT 51.820 59.780 52.050 60.890 ;
        RECT 24.200 53.820 26.200 54.050 ;
        RECT 24.940 52.650 25.240 53.820 ;
        RECT 26.380 52.650 26.680 54.610 ;
        RECT 24.940 52.350 26.680 52.650 ;
        RECT 24.940 48.710 25.240 52.350 ;
        RECT 58.960 51.800 59.320 60.890 ;
        RECT 65.940 60.880 72.550 61.420 ;
        RECT 72.320 59.820 72.550 60.880 ;
        RECT 73.610 61.420 73.840 62.820 ;
        RECT 73.610 61.060 77.060 61.420 ;
        RECT 73.610 59.820 73.840 61.060 ;
        RECT 76.700 51.800 77.060 61.060 ;
        RECT 79.200 56.920 79.590 66.015 ;
        RECT 81.750 61.750 82.770 62.670 ;
        RECT 79.200 56.910 80.180 56.920 ;
        RECT 79.200 56.540 80.225 56.910 ;
        RECT 79.200 56.530 80.180 56.540 ;
        RECT 58.960 51.440 77.060 51.800 ;
        RECT 24.130 48.480 26.130 48.710 ;
        RECT 26.335 48.410 26.565 48.430 ;
        RECT 26.335 47.970 26.690 48.410 ;
        RECT 24.130 47.690 26.130 47.920 ;
        RECT 24.940 45.530 25.200 47.690 ;
        RECT 26.430 45.530 26.690 47.970 ;
        RECT 24.940 45.270 45.150 45.530 ;
        RECT 48.820 45.270 57.360 45.530 ;
        RECT 24.940 42.130 25.200 45.270 ;
        RECT 24.200 41.900 26.200 42.130 ;
        RECT 58.960 35.640 59.320 51.440 ;
        RECT 60.205 45.245 77.715 45.550 ;
        RECT 60.260 45.240 77.715 45.245 ;
        RECT 81.800 38.570 82.720 61.750 ;
        RECT 90.720 56.905 91.065 94.870 ;
        RECT 85.260 56.560 91.065 56.905 ;
        RECT 96.930 86.740 115.350 87.060 ;
        RECT 96.930 45.550 97.250 86.740 ;
        RECT 115.030 85.070 115.350 86.740 ;
        RECT 115.030 84.840 115.395 85.070 ;
        RECT 115.030 84.820 115.350 84.840 ;
        RECT 114.890 80.750 115.120 84.680 ;
        RECT 83.970 45.230 97.250 45.550 ;
        RECT 110.670 80.330 115.120 80.750 ;
        RECT 110.670 44.090 111.090 80.330 ;
        RECT 114.890 79.680 115.120 80.330 ;
        RECT 115.380 81.720 115.610 84.680 ;
        RECT 115.380 80.440 118.650 81.720 ;
        RECT 115.380 79.680 115.610 80.440 ;
        RECT 103.240 43.670 111.090 44.090 ;
        RECT 103.240 38.570 103.660 43.670 ;
        RECT 81.800 37.850 106.830 38.570 ;
        RECT 105.910 37.605 106.830 37.850 ;
        RECT 105.875 36.710 106.870 37.605 ;
        RECT 58.910 35.280 59.370 35.640 ;
        RECT 58.910 31.950 59.370 32.310 ;
        RECT 58.960 31.640 59.320 31.950 ;
        RECT 60.770 31.640 61.000 33.360 ;
        RECT 58.960 31.280 61.000 31.640 ;
        RECT 60.770 29.360 61.000 31.280 ;
        RECT 105.860 29.075 106.870 29.985 ;
        RECT 105.910 27.050 106.820 29.075 ;
        RECT 110.650 27.050 110.880 33.360 ;
        RECT 105.910 26.140 110.880 27.050 ;
        RECT 110.650 17.360 110.880 26.140 ;
      LAYER via ;
        RECT 65.930 69.640 66.470 70.180 ;
        RECT 81.780 69.595 82.730 70.545 ;
        RECT 195.695 109.090 196.105 109.500 ;
        RECT 202.110 109.100 202.510 109.500 ;
        RECT 65.940 63.840 66.480 64.380 ;
        RECT 81.800 61.750 82.720 62.670 ;
        RECT 79.805 56.540 80.175 56.910 ;
        RECT 44.840 45.270 45.100 45.530 ;
        RECT 48.870 45.270 49.130 45.530 ;
        RECT 57.050 45.270 57.310 45.530 ;
        RECT 60.255 45.245 60.560 45.550 ;
        RECT 77.355 45.240 77.665 45.550 ;
        RECT 85.310 56.560 85.655 56.905 ;
        RECT 84.020 45.230 84.340 45.550 ;
        RECT 117.320 80.440 118.600 81.720 ;
        RECT 105.925 36.710 106.820 37.605 ;
        RECT 58.960 35.280 59.320 35.640 ;
        RECT 58.960 31.950 59.320 32.310 ;
        RECT 105.910 29.075 106.820 29.985 ;
      LAYER met2 ;
        RECT 195.695 109.500 196.105 109.550 ;
        RECT 202.110 109.500 202.510 109.550 ;
        RECT 195.695 109.090 202.510 109.500 ;
        RECT 195.695 109.040 196.105 109.090 ;
        RECT 202.110 109.050 202.510 109.090 ;
        RECT 117.320 81.760 118.600 81.770 ;
        RECT 119.310 81.760 120.650 81.800 ;
        RECT 117.300 80.420 120.650 81.760 ;
        RECT 117.320 80.410 120.650 80.420 ;
        RECT 117.320 80.390 118.600 80.410 ;
        RECT 119.310 80.360 120.650 80.410 ;
        RECT 65.930 64.430 66.470 70.230 ;
        RECT 65.930 63.830 66.480 64.430 ;
        RECT 65.940 63.790 66.480 63.830 ;
        RECT 81.780 61.710 82.730 70.595 ;
        RECT 81.800 61.700 82.720 61.710 ;
        RECT 79.805 56.910 80.175 56.960 ;
        RECT 85.310 56.910 85.655 56.955 ;
        RECT 79.805 56.540 85.660 56.910 ;
        RECT 79.805 56.490 80.175 56.540 ;
        RECT 85.310 56.510 85.655 56.540 ;
        RECT 44.840 45.530 45.100 45.580 ;
        RECT 48.870 45.530 49.130 45.580 ;
        RECT 44.840 45.270 49.130 45.530 ;
        RECT 44.840 45.220 45.100 45.270 ;
        RECT 48.870 45.220 49.130 45.270 ;
        RECT 57.050 45.550 57.310 45.580 ;
        RECT 60.255 45.550 60.560 45.600 ;
        RECT 77.355 45.550 77.665 45.600 ;
        RECT 84.020 45.550 84.340 45.600 ;
        RECT 57.050 45.245 60.560 45.550 ;
        RECT 57.050 45.220 57.310 45.245 ;
        RECT 60.255 45.195 60.560 45.245 ;
        RECT 77.350 45.230 84.340 45.550 ;
        RECT 77.355 45.190 77.665 45.230 ;
        RECT 84.020 45.180 84.340 45.230 ;
        RECT 58.960 31.900 59.320 35.690 ;
        RECT 105.925 30.880 106.820 37.655 ;
        RECT 105.910 29.025 106.820 30.880 ;
      LAYER via2 ;
        RECT 119.310 80.410 120.650 81.750 ;
      LAYER met3 ;
        RECT 119.280 81.775 121.380 81.790 ;
        RECT 119.260 81.770 121.380 81.775 ;
        RECT 119.260 80.385 122.740 81.770 ;
        RECT 119.280 80.360 122.740 80.385 ;
      LAYER via3 ;
        RECT 121.280 80.360 122.690 81.770 ;
      LAYER met4 ;
        RECT 132.615 85.715 156.885 115.325 ;
        RECT 160.615 85.715 184.885 115.325 ;
        RECT 141.130 83.180 148.230 85.715 ;
        RECT 169.130 83.180 176.230 85.715 ;
        RECT 141.130 81.840 176.230 83.180 ;
        RECT 122.690 81.800 176.230 81.840 ;
        RECT 121.260 80.360 176.230 81.800 ;
        RECT 121.275 80.355 122.695 80.360 ;
        RECT 141.130 79.040 176.230 80.360 ;
        RECT 141.130 77.325 148.230 79.040 ;
        RECT 169.130 77.325 176.230 79.040 ;
        RECT 132.615 47.715 156.885 77.325 ;
        RECT 160.615 47.715 184.885 77.325 ;
  END
END tt_um_keremergunay_two_stage_opamp
END LIBRARY


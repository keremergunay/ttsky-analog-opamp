magic
tech sky130B
magscale 1 2
timestamp 1768743919
<< metal1 >>
rect 12040 32372 12050 32373
rect 12034 31979 12050 32372
rect 12444 31979 12454 32373
rect 12034 28556 12450 31979
rect 12045 27643 12440 28556
rect 43466 18049 43688 18050
rect 43464 17851 43474 18049
rect 43672 17851 43688 18049
rect 43466 16261 43688 17851
rect 14310 13080 14852 13090
rect 9956 13004 10652 13006
rect 9956 12994 10824 13004
rect 9956 12806 10716 12994
rect 10904 12806 10914 12994
rect 14310 12892 14744 13080
rect 14932 12892 14942 13080
rect 14310 12884 14852 12892
rect 10580 12798 10824 12806
rect 2650 6858 2854 6882
rect 2650 6654 3074 6858
rect 2650 4895 2854 6654
rect 2648 4709 2658 4895
rect 2844 4709 2854 4895
rect 2650 4708 2854 4709
rect 14874 1726 15087 2094
rect 14874 1513 15299 1726
rect 15086 1436 15299 1513
rect 14526 1424 15416 1436
rect 14526 1005 14542 1424
rect 14961 1005 15416 1424
rect 14526 988 15416 1005
<< via1 >>
rect 12050 31979 12444 32373
rect 43474 17851 43672 18049
rect 10716 12806 10904 12994
rect 14744 12892 14932 13080
rect 2658 4709 2844 4895
rect 14542 1005 14961 1424
<< metal2 >>
rect 12050 33000 12446 33010
rect 12050 32608 12054 33000
rect 12050 32598 12446 32608
rect 12050 32373 12444 32598
rect 12050 31969 12444 31979
rect 43482 18388 43670 18396
rect 43474 18386 43672 18388
rect 43474 18198 43482 18386
rect 43670 18198 43672 18386
rect 43474 18049 43672 18198
rect 43474 17841 43672 17851
rect 14744 13082 14932 13090
rect 15008 13082 15192 13084
rect 14744 13080 15194 13082
rect 10716 12996 10904 13004
rect 10980 12996 11164 12998
rect 10716 12994 11166 12996
rect 10904 12988 11166 12994
rect 10904 12806 10980 12988
rect 10716 12804 10980 12806
rect 11164 12804 11166 12988
rect 14932 13074 15194 13080
rect 14932 12892 15008 13074
rect 14744 12890 15008 12892
rect 15192 12890 15194 13074
rect 14744 12882 14932 12890
rect 15008 12880 15192 12890
rect 10716 12796 10904 12804
rect 10980 12794 11164 12804
rect 2658 4895 2844 4905
rect 2654 4709 2658 4732
rect 2654 4556 2844 4709
rect 2654 4546 2846 4556
rect 2654 4358 2658 4546
rect 2654 4356 2846 4358
rect 2658 4348 2846 4356
rect 14542 1424 14961 1434
rect 14125 1416 14542 1424
rect 13720 1406 14542 1416
rect 14136 1006 14542 1406
rect 14136 990 14150 1006
rect 14536 1005 14542 1006
rect 14542 995 14961 1005
rect 13720 988 14150 990
rect 13720 980 14136 988
<< via2 >>
rect 12054 32608 12446 33000
rect 43482 18198 43670 18386
rect 10980 12804 11164 12988
rect 15008 12890 15192 13074
rect 2658 4358 2846 4546
rect 13720 990 14136 1406
<< metal3 >>
rect 12054 33738 12446 33746
rect 12046 33338 12056 33738
rect 12456 33338 12466 33738
rect 12054 33005 12446 33338
rect 12044 33000 12456 33005
rect 12044 32608 12054 33000
rect 12446 32608 12456 33000
rect 12044 32603 12456 32608
rect 43482 18702 43670 18704
rect 43474 18522 43484 18702
rect 43664 18522 43674 18702
rect 43482 18391 43670 18522
rect 43472 18386 43680 18391
rect 43472 18198 43482 18386
rect 43670 18198 43680 18386
rect 43472 18193 43680 18198
rect 14998 13074 15202 13079
rect 10970 12988 11174 12993
rect 10970 12804 10980 12988
rect 11164 12808 11276 12988
rect 11456 12808 11466 12988
rect 14998 12890 15008 13074
rect 15192 12894 15304 13074
rect 15484 12894 15494 13074
rect 15192 12890 15484 12894
rect 14998 12885 15202 12890
rect 11164 12804 11456 12808
rect 10970 12799 11174 12804
rect 2648 4546 2856 4551
rect 2648 4358 2658 4546
rect 2846 4358 2856 4546
rect 2648 4353 2856 4358
rect 2658 4234 2846 4353
rect 2644 4054 2654 4234
rect 2834 4054 2846 4234
rect 2658 4046 2846 4054
rect 13710 1406 14146 1411
rect 13020 1398 13720 1406
rect 13020 998 13040 1398
rect 13440 998 13720 1398
rect 13020 990 13720 998
rect 14136 990 14146 1406
rect 13020 985 14146 990
rect 13020 976 13856 985
<< via3 >>
rect 12056 33338 12456 33738
rect 43484 18522 43664 18702
rect 11276 12808 11456 12988
rect 15304 12894 15484 13074
rect 2654 4054 2834 4234
rect 13040 998 13440 1398
<< metal4 >>
rect 5934 44950 5994 45150
rect 6486 44950 6546 45150
rect 7038 44950 7098 45150
rect 7590 44950 7650 45150
rect 8142 44950 8202 45150
rect 8694 44950 8754 45150
rect 9246 44950 9306 45150
rect 9798 44950 9858 45150
rect 10350 44950 10410 45150
rect 10902 44950 10962 45150
rect 11454 44950 11514 45150
rect 12006 44950 12066 45150
rect 12558 44950 12618 45150
rect 13110 44950 13170 45150
rect 13662 44950 13722 45150
rect 14214 44950 14274 45150
rect 14766 44950 14826 45150
rect 15318 44950 15378 45150
rect 15870 44950 15930 45150
rect 16422 44950 16482 45150
rect 16974 44950 17034 45150
rect 17526 44950 17586 45150
rect 18078 44950 18138 45150
rect 18630 44950 18690 45150
rect 19182 44950 19242 45150
rect 19734 44950 19794 45150
rect 20286 44950 20346 45150
rect 20838 44950 20898 45150
rect 21390 44950 21450 45150
rect 21942 44950 22002 45150
rect 22494 44950 22554 45150
rect 23046 44950 23106 45150
rect 23598 44950 23658 45150
rect 24150 44950 24210 45150
rect 24702 44950 24762 45150
rect 25254 44950 25314 45150
rect 25806 44950 25866 45150
rect 26358 44950 26418 45150
rect 26910 44950 26970 45150
rect 27462 44950 27522 45150
rect 28014 44950 28074 45150
rect 28566 44950 28626 45150
rect 29118 44950 29178 45150
rect 0 44382 4586 44782
rect 0 998 400 44382
rect 600 1398 1000 44150
rect 4186 34592 4586 44382
rect 4186 34192 12456 34592
rect 12056 33739 12456 34192
rect 12055 33738 12457 33739
rect 12055 33338 12056 33738
rect 12456 33338 12457 33738
rect 12055 33337 12457 33338
rect 6600 26992 40428 27172
rect 6600 8520 6780 26992
rect 40248 23052 40428 26992
rect 40248 22872 40844 23052
rect 40664 18702 40844 22872
rect 43483 18702 43665 18703
rect 40664 18522 43484 18702
rect 43664 18522 43665 18702
rect 43483 18521 43665 18522
rect 15303 13074 15485 13075
rect 11446 12989 12576 12998
rect 11275 12988 12576 12989
rect 11275 12808 11276 12988
rect 11456 12818 12576 12988
rect 15303 12894 15304 13074
rect 15484 12894 25046 13074
rect 15303 12893 15485 12894
rect 11456 12808 11570 12818
rect 11275 12807 11457 12808
rect 12396 11058 12576 12818
rect 12396 10878 23738 11058
rect 6600 8340 17424 8520
rect 2653 4234 2835 4235
rect 2653 4054 2654 4234
rect 2834 4054 2835 4234
rect 2653 4053 2835 4054
rect 2654 3990 2834 4053
rect 2654 3810 16566 3990
rect 13039 1398 13441 1399
rect 600 998 13040 1398
rect 13440 998 13441 1398
rect 13039 997 13441 998
rect 16386 666 16566 3810
rect 17244 2550 17424 8340
rect 23558 7908 23738 10878
rect 24866 8678 25046 12894
rect 24866 8498 30342 8678
rect 23558 7728 26478 7908
rect 17244 2370 22614 2550
rect 16386 486 18750 666
rect 3114 -2 3294 198
rect 6978 -2 7158 198
rect 10842 -2 11022 198
rect 14706 -2 14886 198
rect 18570 -2 18750 486
rect 22434 -2 22614 2370
rect 26298 -2 26478 7728
rect 30162 -2 30342 8498
use two_stage_opamp  two_stage_opamp_0 ~/Desktop/design/mag/Final_Project
timestamp 1768091639
transform 1 0 -308 0 1 11032
box 3266 -9126 44228 16662
<< labels >>
flabel metal4 s 28566 44950 28626 45150 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29118 44950 29178 45150 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28014 44950 28074 45150 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30162 -2 30342 198 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26298 -2 26478 198 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22434 -2 22614 198 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18570 -2 18750 198 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14706 -2 14886 198 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 10842 -2 11022 198 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 6978 -2 7158 198 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3114 -2 3294 198 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27462 44950 27522 45150 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 26910 44950 26970 45150 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26358 44950 26418 45150 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 25806 44950 25866 45150 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25254 44950 25314 45150 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24702 44950 24762 45150 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24150 44950 24210 45150 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23598 44950 23658 45150 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23046 44950 23106 45150 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22494 44950 22554 45150 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 21942 44950 22002 45150 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21390 44950 21450 45150 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20838 44950 20898 45150 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20286 44950 20346 45150 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19734 44950 19794 45150 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19182 44950 19242 45150 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9798 44950 9858 45150 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 9246 44950 9306 45150 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 8694 44950 8754 45150 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 8142 44950 8202 45150 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 7590 44950 7650 45150 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 7038 44950 7098 45150 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 6486 44950 6546 45150 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 5934 44950 5994 45150 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 14214 44950 14274 45150 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 13662 44950 13722 45150 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 13110 44950 13170 45150 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 12558 44950 12618 45150 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 12006 44950 12066 45150 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 11454 44950 11514 45150 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 10902 44950 10962 45150 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 10350 44950 10410 45150 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 18630 44950 18690 45150 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 18078 44950 18138 45150 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 17526 44950 17586 45150 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 16974 44950 17034 45150 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 16422 44950 16482 45150 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 15870 44950 15930 45150 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 15318 44950 15378 45150 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 14766 44950 14826 45150 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 0 998 400 44150 1 FreeSans 2 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 600 998 1000 44150 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< end >>
